netcdf lon.0.625x0.5 {
dimensions:
	lon = 576 ;

variables:
	float lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;

// global attributes:
		:Conventions = "COARDS" ;
		:Source = "Unknown" ;
		:Title = "Unknown" ;
		:Contact = "Unknown" ;
		:History = "Mon Mar  7 12:42:46 2016: ncks -v lon MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.nc lon.1x1.25.nc\n",
    "Wed Sep 15 22:23:40 2010: ncrename -d record,time /home/mrdamon/ProcessMerra300/MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.nc\n",
    "Mon Sep 13 18:28:53 2010: ncks -v FRLAKE,FRLAND,FRLANDICE,FROCEAN MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.nc 1x1.25.nc\n",
    "Mon Sep 13 18:00:38 2010: ncks -v lev /discover/nobackup/mrdamon/Devel/GmiAutomation/GEOS5DAS-discover/levs.nc --append MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.nc\n",
    "Mon Sep 13 17:57:31 2010: ncwa -a time reduced.1x1.25.nc MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.nc\n",
    "Mon Sep 13 17:56:36 2010: ncks -v FRLAKE,FRLAND,FRLANDICE,FROCEAN MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.nc reduced.1x1.25.nc\n",
    "Mon Sep 13 17:15:43 2010: ncecat MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.1.nc MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.2.nc MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.3.nc MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.4.nc MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.5.nc MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.6.nc MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.8.nc MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.7.nc test.nc\n",
    "Sun Sep 12 17:34:49 2010: ncatted -O -a Met_Data_Name,global,o,c,GMAO_GEOS5MERRA300_1x1%25x72 MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.nc\n",
    "Sun Sep 12 17:34:30 2010: ncatted -O -a Met_Data_Name,global,a,c,GMAO_GEOS5MERRA300_1x1%25x72 MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.nc\n",
    "Thu Sep  9 14:43:04 2010: ncks -v lev /archive/anon/pub/gmidata2/input/metfields/geos5das-merra/1x1.25/2003/MERRA300.prod.assim.20030128.1x1.25.nc --append MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.ncks.nc\n",
    "Thu Sep  9 14:33:55 2010: ncks -v FRLAKE,FRLAND,FRLANDICE,FROCEAN,lon,lat,time MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.nc MERRA300.prod.assim.const_2d_asm_Nx.00000000.1x1.25.ncks.nc\n",
    "File written by GFIO v1.0.8" ;
		:ptop = 0.f ;
		:pint = 0.f ;
		:ks = -1.f ;
		:ak = 0.f ;
		:bk = 0.f ;
		:Met_Data_Name = "GMAO_GEOS5MERRA2_0%625x0%5x72" ;
		:nco_openmp_thread_number = 1 ;
		:NCO = "4.2.3" ;

data:

 lon = 0 , 0.625 , 1.25 , 1.875 , 2.5 , 3.125 , 3.75 , 4.375 , 5 , 5.625 , 
    6.25 , 6.875 , 7.5 , 8.125 , 8.75 , 9.375 , 10 , 10.625 , 11.25 , 
    11.875 , 12.5 , 13.125 , 13.75 , 14.375 , 15 , 15.625 , 16.25 , 16.875 , 
    17.5 , 18.125 , 18.75 , 19.375 , 20 , 20.625 , 21.25 , 21.875 , 22.5 , 
    23.125 , 23.75 , 24.375 , 25 , 25.625 , 26.25 , 26.875 , 27.5 , 28.125 , 
    28.75 , 29.375 , 30 , 30.625 , 31.25 , 31.875 , 32.5 , 33.125 , 33.75 , 
    34.375 , 35 , 35.625 , 36.25 , 36.875 , 37.5 , 38.125 , 38.75 , 39.375 , 
    40 , 40.625 , 41.25 , 41.875 , 42.5 , 43.125 , 43.75 , 44.375 , 45 , 
    45.625 , 46.25 , 46.875 , 47.5 , 48.125 , 48.75 , 49.375 , 50 , 50.625 , 
    51.25 , 51.875 , 52.5 , 53.125 , 53.75 , 54.375 , 55 , 55.625 , 56.25 , 
    56.875 , 57.5 , 58.125 , 58.75 , 59.375 , 60 , 60.625 , 61.25 , 61.875 , 
    62.5 , 63.125 , 63.75 , 64.375 , 65 , 65.625 , 66.25 , 66.875 , 67.5 , 
    68.125 , 68.75 , 69.375 , 70 , 70.625 , 71.25 , 71.875 , 72.5 , 73.125 , 
    73.75 , 74.375 , 75 , 75.625 , 76.25 , 76.875 , 77.5 , 78.125 , 78.75 , 
    79.375 , 80 , 80.625 , 81.25 , 81.875 , 82.5 , 83.125 , 83.75 , 84.375 , 
    85 , 85.625 , 86.25 , 86.875 , 87.5 , 88.125 , 88.75 , 89.375 , 90 , 
    90.625 , 91.25 , 91.875 , 92.5 , 93.125 , 93.75 , 94.375 , 95 , 95.625 , 
    96.25 , 96.875 , 97.5 , 98.125 , 98.75 , 99.375 , 100 , 100.625 , 
    101.25 , 101.875 , 102.5 , 103.125 , 103.75 , 104.375 , 105 , 105.625 , 
    106.25 , 106.875 , 107.5 , 108.125 , 108.75 , 109.375 , 110 , 110.625 , 
    111.25 , 111.875 , 112.5 , 113.125 , 113.75 , 114.375 , 115 , 115.625 , 
    116.25 , 116.875 , 117.5 , 118.125 , 118.75 , 119.375 , 120 , 120.625 , 
    121.25 , 121.875 , 122.5 , 123.125 , 123.75 , 124.375 , 125 , 125.625 , 
    126.25 , 126.875 , 127.5 , 128.125 , 128.75 , 129.375 , 130 , 130.625 , 
    131.25 , 131.875 , 132.5 , 133.125 , 133.75 , 134.375 , 135 , 135.625 , 
    136.25 , 136.875 , 137.5 , 138.125 , 138.75 , 139.375 , 140 , 140.625 , 
    141.25 , 141.875 , 142.5 , 143.125 , 143.75 , 144.375 , 145 , 145.625 , 
    146.25 , 146.875 , 147.5 , 148.125 , 148.75 , 149.375 , 150 , 150.625 , 
    151.25 , 151.875 , 152.5 , 153.125 , 153.75 , 154.375 , 155 , 155.625 , 
    156.25 , 156.875 , 157.5 , 158.125 , 158.75 , 159.375 , 160 , 160.625 , 
    161.25 , 161.875 , 162.5 , 163.125 , 163.75 , 164.375 , 165 , 165.625 , 
    166.25 , 166.875 , 167.5 , 168.125 , 168.75 , 169.375 , 170 , 170.625 , 
    171.25 , 171.875 , 172.5 , 173.125 , 173.75 , 174.375 , 175 , 175.625 , 
    176.25 , 176.875 , 177.5 , 178.125 , 178.75 , 179.375 , 180 , 180.625 , 
    181.25 , 181.875 , 182.5 , 183.125 , 183.75 , 184.375 , 185 , 185.625 , 
    186.25 , 186.875 , 187.5 , 188.125 , 188.75 , 189.375 , 190 , 190.625 , 
    191.25 , 191.875 , 192.5 , 193.125 , 193.75 , 194.375 , 195 , 195.625 , 
    196.25 , 196.875 , 197.5 , 198.125 , 198.75 , 199.375 , 200 , 200.625 , 
    201.25 , 201.875 , 202.5 , 203.125 , 203.75 , 204.375 , 205 , 205.625 , 
    206.25 , 206.875 , 207.5 , 208.125 , 208.75 , 209.375 , 210 , 210.625 , 
    211.25 , 211.875 , 212.5 , 213.125 , 213.75 , 214.375 , 215 , 215.625 , 
    216.25 , 216.875 , 217.5 , 218.125 , 218.75 , 219.375 , 220 , 220.625 , 
    221.25 , 221.875 , 222.5 , 223.125 , 223.75 , 224.375 , 225 , 225.625 , 
    226.25 , 226.875 , 227.5 , 228.125 , 228.75 , 229.375 , 230 , 230.625 , 
    231.25 , 231.875 , 232.5 , 233.125 , 233.75 , 234.375 , 235 , 235.625 , 
    236.25 , 236.875 , 237.5 , 238.125 , 238.75 , 239.375 , 240 , 240.625 , 
    241.25 , 241.875 , 242.5 , 243.125 , 243.75 , 244.375 , 245 , 245.625 , 
    246.25 , 246.875 , 247.5 , 248.125 , 248.75 , 249.375 , 250 , 250.625 , 
    251.25 , 251.875 , 252.5 , 253.125 , 253.75 , 254.375 , 255 , 255.625 , 
    256.25 , 256.875 , 257.5 , 258.125 , 258.75 , 259.375 , 260 , 260.625 , 
    261.25 , 261.875 , 262.5 , 263.125 , 263.75 , 264.375 , 265 , 265.625 , 
    266.25 , 266.875 , 267.5 , 268.125 , 268.75 , 269.375 , 270 , 270.625 , 
    271.25 , 271.875 , 272.5 , 273.125 , 273.75 , 274.375 , 275 , 275.625 , 
    276.25 , 276.875 , 277.5 , 278.125 , 278.75 , 279.375 , 280 , 280.625 , 
    281.25 , 281.875 , 282.5 , 283.125 , 283.75 , 284.375 , 285 , 285.625 , 
    286.25 , 286.875 , 287.5 , 288.125 , 288.75 , 289.375 , 290 , 290.625 , 
    291.25 , 291.875 , 292.5 , 293.125 , 293.75 , 294.375 , 295 , 295.625 , 
    296.25 , 296.875 , 297.5 , 298.125 , 298.75 , 299.375 , 300 , 300.625 , 
    301.25 , 301.875 , 302.5 , 303.125 , 303.75 , 304.375 , 305 , 305.625 , 
    306.25 , 306.875 , 307.5 , 308.125 , 308.75 , 309.375 , 310 , 310.625 , 
    311.25 , 311.875 , 312.5 , 313.125 , 313.75 , 314.375 , 315 , 315.625 , 
    316.25 , 316.875 , 317.5 , 318.125 , 318.75 , 319.375 , 320 , 320.625 , 
    321.25 , 321.875 , 322.5 , 323.125 , 323.75 , 324.375 , 325 , 325.625 , 
    326.25 , 326.875 , 327.5 , 328.125 , 328.75 , 329.375 , 330 , 330.625 , 
    331.25 , 331.875 , 332.5 , 333.125 , 333.75 , 334.375 , 335 , 335.625 , 
    336.25 , 336.875 , 337.5 , 338.125 , 338.75 , 339.375 , 340 , 340.625 , 
    341.25 , 341.875 , 342.5 , 343.125 , 343.75 , 344.375 , 345 , 345.625 , 
    346.25 , 346.875 , 347.5 , 348.125 , 348.75 , 349.375 , 350 , 350.625 , 
    351.25 , 351.875 , 352.5 , 353.125 , 353.75 , 354.375 , 355 , 355.625 , 
    356.25 , 356.875 , 357.5 , 358.125 , 358.75 , 359.375  ;
}
