netcdf lon.1x1.25 {
dimensions:
	lon = 288 ;

variables:
	float lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;

// global attributes:
		:Conventions = "COARDS" ;
		:Source = "Unknown" ;
		:Title = "Unknown" ;
		:Contact = "Unknown" ;

data:

 lon = 0 , 1.25 , 2.5 , 3.75 , 5 , 6.25 , 7.5 , 8.75 , 10 , 11.25 , 12.5 , 
    13.75 , 15 , 16.25 , 17.5 , 18.75 , 20 , 21.25 , 22.5 , 23.75 , 25 , 
    26.25 , 27.5 , 28.75 , 30 , 31.25 , 32.5 , 33.75 , 35 , 36.25 , 37.5 , 
    38.75 , 40 , 41.25 , 42.5 , 43.75 , 45 , 46.25 , 47.5 , 48.75 , 50 , 
    51.25 , 52.5 , 53.75 , 55 , 56.25 , 57.5 , 58.75 , 60 , 61.25 , 62.5 , 
    63.75 , 65 , 66.25 , 67.5 , 68.75 , 70 , 71.25 , 72.5 , 73.75 , 75 , 
    76.25 , 77.5 , 78.75 , 80 , 81.25 , 82.5 , 83.75 , 85 , 86.25 , 87.5 , 
    88.75 , 90 , 91.25 , 92.5 , 93.75 , 95 , 96.25 , 97.5 , 98.75 , 100 , 
    101.25 , 102.5 , 103.75 , 105 , 106.25 , 107.5 , 108.75 , 110 , 111.25 , 
    112.5 , 113.75 , 115 , 116.25 , 117.5 , 118.75 , 120 , 121.25 , 122.5 , 
    123.75 , 125 , 126.25 , 127.5 , 128.75 , 130 , 131.25 , 132.5 , 133.75 , 
    135 , 136.25 , 137.5 , 138.75 , 140 , 141.25 , 142.5 , 143.75 , 145 , 
    146.25 , 147.5 , 148.75 , 150 , 151.25 , 152.5 , 153.75 , 155 , 156.25 , 
    157.5 , 158.75 , 160 , 161.25 , 162.5 , 163.75 , 165 , 166.25 , 167.5 , 
    168.75 , 170 , 171.25 , 172.5 , 173.75 , 175 , 176.25 , 177.5 , 178.75 , 
    180 , 181.25 , 182.5 , 183.75 , 185 , 186.25 , 187.5 , 188.75 , 190 , 
    191.25 , 192.5 , 193.75 , 195 , 196.25 , 197.5 , 198.75 , 200 , 201.25 , 
    202.5 , 203.75 , 205 , 206.25 , 207.5 , 208.75 , 210 , 211.25 , 212.5 , 
    213.75 , 215 , 216.25 , 217.5 , 218.75 , 220 , 221.25 , 222.5 , 223.75 , 
    225 , 226.25 , 227.5 , 228.75 , 230 , 231.25 , 232.5 , 233.75 , 235 , 
    236.25 , 237.5 , 238.75 , 240 , 241.25 , 242.5 , 243.75 , 245 , 246.25 , 
    247.5 , 248.75 , 250 , 251.25 , 252.5 , 253.75 , 255 , 256.25 , 257.5 , 
    258.75 , 260 , 261.25 , 262.5 , 263.75 , 265 , 266.25 , 267.5 , 268.75 , 
    270 , 271.25 , 272.5 , 273.75 , 275 , 276.25 , 277.5 , 278.75 , 280 , 
    281.25 , 282.5 , 283.75 , 285 , 286.25 , 287.5 , 288.75 , 290 , 291.25 , 
    292.5 , 293.75 , 295 , 296.25 , 297.5 , 298.75 , 300 , 301.25 , 302.5 , 
    303.75 , 305 , 306.25 , 307.5 , 308.75 , 310 , 311.25 , 312.5 , 313.75 , 
    315 , 316.25 , 317.5 , 318.75 , 320 , 321.25 , 322.5 , 323.75 , 325 , 
    326.25 , 327.5 , 328.75 , 330 , 331.25 , 332.5 , 333.75 , 335 , 336.25 , 
    337.5 , 338.75 , 340 , 341.25 , 342.5 , 343.75 , 345 , 346.25 , 347.5 , 
    348.75 , 350 , 351.25 , 352.5 , 353.75 , 355 , 356.25 , 357.5 , 358.75  ;
}
