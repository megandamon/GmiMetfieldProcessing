netcdf lon.2x2.5 {
dimensions:
	lon = 144 ;

variables:
	float lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;

// global attributes:
		:Conventions = "COARDS" ;
		:Source = "Unknown" ;
		:Title = "Unknown" ;
		:Contact = "Unknown" ;
		:History = "Mon Mar  7 12:43:00 2016: ncks -v lon MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.nc lon.2x2.5.nc\n",
    "Wed Sep 15 18:12:59 2010: ncrename -v time,time1 /home/mrdamon/ProcessMerra300/MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.nc\n",
    "Mon Sep 13 18:29:03 2010: ncks -v FRLAKE,FRLAND,FRLANDICE,FROCEAN MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.nc 2x2.5.nc\n",
    "Mon Sep 13 18:23:40 2010: ncrename -v am,am3 -v bm,bm3 MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.nc\n",
    "Mon Sep 13 18:17:25 2010: ncrename -v am,am_2 -v bm,bm_2 MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.nc\n",
    "Mon Sep 13 18:16:41 2010: ncrename -v lev72,lev MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.nc\n",
    "Mon Sep 13 18:14:29 2010: ncrename -v lev,lev72 MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.nc\n",
    "Mon Sep 13 18:00:35 2010: ncks -v lev /discover/nobackup/mrdamon/Devel/GmiAutomation/GEOS5DAS-discover/levs.nc --append MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.nc\n",
    "Mon Sep 13 17:56:26 2010: ncks -v FRLAKE,FRLAND,FRLANDICE,FROCEAN MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.nc reduced.2x2.5.nc\n",
    "Mon Sep 13 17:55:23 2010: ncrename -d record,time MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.nc\n",
    "Mon Sep 13 17:53:52 2010: ncwa -a time test.nc MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.removed.nc\n",
    "Mon Sep 13 17:53:05 2010: ncecat MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.1.nc MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.2.nc MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.4.nc MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.3.nc MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.6.nc MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.5.nc MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.7.nc MERRA300.prod.assim.const_2d_asm_Nx.00000000.2x2.5.8.nc test.nc\n",
    "File written by GFIO v1.0.8" ;
		:ptop = 0.f ;
		:pint = 0.f ;
		:ks = -1.f ;
		:ak = 0.f ;
		:bk = 0.f ;
		:nco_openmp_thread_number = 1 ;
		:Met_Data_Name = "GMAO_GEOS5MERRA2_2x2%5x72" ;
		:NCO = "4.2.3" ;

data:

 lon = 0 , 2.5 , 5 , 7.5 , 10 , 12.5 , 15 , 17.5 , 20 , 22.5 , 25 , 27.5 , 
    30 , 32.5 , 35 , 37.5 , 40 , 42.5 , 45 , 47.5 , 50 , 52.5 , 55 , 57.5 , 
    60 , 62.5 , 65 , 67.5 , 70 , 72.5 , 75 , 77.5 , 80 , 82.5 , 85 , 87.5 , 
    90 , 92.5 , 95 , 97.5 , 100 , 102.5 , 105 , 107.5 , 110 , 112.5 , 115 , 
    117.5 , 120 , 122.5 , 125 , 127.5 , 130 , 132.5 , 135 , 137.5 , 140 , 
    142.5 , 145 , 147.5 , 150 , 152.5 , 155 , 157.5 , 160 , 162.5 , 165 , 
    167.5 , 170 , 172.5 , 175 , 177.5 , 180 , 182.5 , 185 , 187.5 , 190 , 
    192.5 , 195 , 197.5 , 200 , 202.5 , 205 , 207.5 , 210 , 212.5 , 215 , 
    217.5 , 220 , 222.5 , 225 , 227.5 , 230 , 232.5 , 235 , 237.5 , 240 , 
    242.5 , 245 , 247.5 , 250 , 252.5 , 255 , 257.5 , 260 , 262.5 , 265 , 
    267.5 , 270 , 272.5 , 275 , 277.5 , 280 , 282.5 , 285 , 287.5 , 290 , 
    292.5 , 295 , 297.5 , 300 , 302.5 , 305 , 307.5 , 310 , 312.5 , 315 , 
    317.5 , 320 , 322.5 , 325 , 327.5 , 330 , 332.5 , 335 , 337.5 , 340 , 
    342.5 , 345 , 347.5 , 350 , 352.5 , 355 , 357.5  ;
}
